`default_nettype none

module aludec();
endmodule

`default_nettype wire
