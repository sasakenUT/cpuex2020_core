`default_nettype none

module datapath();
endmodule

`default_nettype wire
