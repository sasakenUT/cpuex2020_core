`default_nettype none

module riscv();
endmodule

`default_nettype wire
