`default_nettype none

module controller();
endmodule

`default_nettype wire
